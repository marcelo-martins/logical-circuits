LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY UC IS 
		PORT (
			--io
		);
END ENTITY;

architecture fulltrab of UC is

--ESTADOS DA MAQUINA DE CAFFERSON
type estado_maq is (escolhendo_cafe, pagando, troco, fazendo_cafe);




begin




end fulltrab
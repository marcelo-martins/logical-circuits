LIBRARY ieee;
USE ieee.std_logic_1164.ALL;


ENTITY bico_cafe IS 
		PORT (
			dispence_coffee		: IN 	STD_LOGIC; 
			dispensing_coffee	   : OUT	STD_LOGIC;
		);
END ENTITY;

